##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Tue Apr 20 01:22:18 2021
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ensc450
  CLASS BLOCK ;
  SIZE 649.990000 BY 650.020000 ;
  FOREIGN ensc450 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
  END clk
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 191.770000 649.950000 191.840000 650.020000 ;
    END
  END resetn
  PIN EXT_NREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 436.835000 0.070000 436.905000 ;
    END
  END EXT_NREADY
  PIN EXT_BUSY
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 199.370000 649.950000 199.440000 650.020000 ;
    END
  END EXT_BUSY
  PIN EXT_MR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 206.970000 649.950000 207.040000 650.020000 ;
    END
  END EXT_MR
  PIN EXT_MW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 214.570000 649.950000 214.640000 650.020000 ;
    END
  END EXT_MW
  PIN EXT_ADDRBUS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 222.170000 649.950000 222.240000 650.020000 ;
    END
  END EXT_ADDRBUS[31]
  PIN EXT_ADDRBUS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 229.770000 649.950000 229.840000 650.020000 ;
    END
  END EXT_ADDRBUS[30]
  PIN EXT_ADDRBUS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 237.370000 649.950000 237.440000 650.020000 ;
    END
  END EXT_ADDRBUS[29]
  PIN EXT_ADDRBUS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 244.970000 649.950000 245.040000 650.020000 ;
    END
  END EXT_ADDRBUS[28]
  PIN EXT_ADDRBUS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 252.570000 649.950000 252.640000 650.020000 ;
    END
  END EXT_ADDRBUS[27]
  PIN EXT_ADDRBUS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 260.170000 649.950000 260.240000 650.020000 ;
    END
  END EXT_ADDRBUS[26]
  PIN EXT_ADDRBUS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 267.770000 649.950000 267.840000 650.020000 ;
    END
  END EXT_ADDRBUS[25]
  PIN EXT_ADDRBUS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 275.370000 649.950000 275.440000 650.020000 ;
    END
  END EXT_ADDRBUS[24]
  PIN EXT_ADDRBUS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 282.970000 649.950000 283.040000 650.020000 ;
    END
  END EXT_ADDRBUS[23]
  PIN EXT_ADDRBUS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 290.570000 649.950000 290.640000 650.020000 ;
    END
  END EXT_ADDRBUS[22]
  PIN EXT_ADDRBUS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 298.170000 649.950000 298.240000 650.020000 ;
    END
  END EXT_ADDRBUS[21]
  PIN EXT_ADDRBUS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 305.770000 649.950000 305.840000 650.020000 ;
    END
  END EXT_ADDRBUS[20]
  PIN EXT_ADDRBUS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 313.370000 649.950000 313.440000 650.020000 ;
    END
  END EXT_ADDRBUS[19]
  PIN EXT_ADDRBUS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 320.970000 649.950000 321.040000 650.020000 ;
    END
  END EXT_ADDRBUS[18]
  PIN EXT_ADDRBUS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 328.570000 649.950000 328.640000 650.020000 ;
    END
  END EXT_ADDRBUS[17]
  PIN EXT_ADDRBUS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 336.170000 649.950000 336.240000 650.020000 ;
    END
  END EXT_ADDRBUS[16]
  PIN EXT_ADDRBUS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 343.770000 649.950000 343.840000 650.020000 ;
    END
  END EXT_ADDRBUS[15]
  PIN EXT_ADDRBUS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 351.370000 649.950000 351.440000 650.020000 ;
    END
  END EXT_ADDRBUS[14]
  PIN EXT_ADDRBUS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 358.970000 649.950000 359.040000 650.020000 ;
    END
  END EXT_ADDRBUS[13]
  PIN EXT_ADDRBUS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 366.570000 649.950000 366.640000 650.020000 ;
    END
  END EXT_ADDRBUS[12]
  PIN EXT_ADDRBUS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.170000 649.950000 374.240000 650.020000 ;
    END
  END EXT_ADDRBUS[11]
  PIN EXT_ADDRBUS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 381.770000 649.950000 381.840000 650.020000 ;
    END
  END EXT_ADDRBUS[10]
  PIN EXT_ADDRBUS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 389.370000 649.950000 389.440000 650.020000 ;
    END
  END EXT_ADDRBUS[9]
  PIN EXT_ADDRBUS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 396.970000 649.950000 397.040000 650.020000 ;
    END
  END EXT_ADDRBUS[8]
  PIN EXT_ADDRBUS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 404.570000 649.950000 404.640000 650.020000 ;
    END
  END EXT_ADDRBUS[7]
  PIN EXT_ADDRBUS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 412.170000 649.950000 412.240000 650.020000 ;
    END
  END EXT_ADDRBUS[6]
  PIN EXT_ADDRBUS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 419.770000 649.950000 419.840000 650.020000 ;
    END
  END EXT_ADDRBUS[5]
  PIN EXT_ADDRBUS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 427.370000 649.950000 427.440000 650.020000 ;
    END
  END EXT_ADDRBUS[4]
  PIN EXT_ADDRBUS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 434.970000 649.950000 435.040000 650.020000 ;
    END
  END EXT_ADDRBUS[3]
  PIN EXT_ADDRBUS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 442.570000 649.950000 442.640000 650.020000 ;
    END
  END EXT_ADDRBUS[2]
  PIN EXT_ADDRBUS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 450.170000 649.950000 450.240000 650.020000 ;
    END
  END EXT_ADDRBUS[1]
  PIN EXT_ADDRBUS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 457.770000 649.950000 457.840000 650.020000 ;
    END
  END EXT_ADDRBUS[0]
  PIN EXT_RDATABUS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 212.835000 0.070000 212.905000 ;
    END
  END EXT_RDATABUS[31]
  PIN EXT_RDATABUS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 219.835000 0.070000 219.905000 ;
    END
  END EXT_RDATABUS[30]
  PIN EXT_RDATABUS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 226.835000 0.070000 226.905000 ;
    END
  END EXT_RDATABUS[29]
  PIN EXT_RDATABUS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 233.835000 0.070000 233.905000 ;
    END
  END EXT_RDATABUS[28]
  PIN EXT_RDATABUS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 240.835000 0.070000 240.905000 ;
    END
  END EXT_RDATABUS[27]
  PIN EXT_RDATABUS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 247.835000 0.070000 247.905000 ;
    END
  END EXT_RDATABUS[26]
  PIN EXT_RDATABUS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 254.835000 0.070000 254.905000 ;
    END
  END EXT_RDATABUS[25]
  PIN EXT_RDATABUS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 261.835000 0.070000 261.905000 ;
    END
  END EXT_RDATABUS[24]
  PIN EXT_RDATABUS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 268.835000 0.070000 268.905000 ;
    END
  END EXT_RDATABUS[23]
  PIN EXT_RDATABUS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 275.835000 0.070000 275.905000 ;
    END
  END EXT_RDATABUS[22]
  PIN EXT_RDATABUS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 282.835000 0.070000 282.905000 ;
    END
  END EXT_RDATABUS[21]
  PIN EXT_RDATABUS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 289.835000 0.070000 289.905000 ;
    END
  END EXT_RDATABUS[20]
  PIN EXT_RDATABUS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 296.835000 0.070000 296.905000 ;
    END
  END EXT_RDATABUS[19]
  PIN EXT_RDATABUS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 303.835000 0.070000 303.905000 ;
    END
  END EXT_RDATABUS[18]
  PIN EXT_RDATABUS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 310.835000 0.070000 310.905000 ;
    END
  END EXT_RDATABUS[17]
  PIN EXT_RDATABUS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 317.835000 0.070000 317.905000 ;
    END
  END EXT_RDATABUS[16]
  PIN EXT_RDATABUS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 324.835000 0.070000 324.905000 ;
    END
  END EXT_RDATABUS[15]
  PIN EXT_RDATABUS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 331.835000 0.070000 331.905000 ;
    END
  END EXT_RDATABUS[14]
  PIN EXT_RDATABUS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 338.835000 0.070000 338.905000 ;
    END
  END EXT_RDATABUS[13]
  PIN EXT_RDATABUS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 345.835000 0.070000 345.905000 ;
    END
  END EXT_RDATABUS[12]
  PIN EXT_RDATABUS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 352.835000 0.070000 352.905000 ;
    END
  END EXT_RDATABUS[11]
  PIN EXT_RDATABUS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 359.835000 0.070000 359.905000 ;
    END
  END EXT_RDATABUS[10]
  PIN EXT_RDATABUS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 366.835000 0.070000 366.905000 ;
    END
  END EXT_RDATABUS[9]
  PIN EXT_RDATABUS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 373.835000 0.070000 373.905000 ;
    END
  END EXT_RDATABUS[8]
  PIN EXT_RDATABUS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 380.835000 0.070000 380.905000 ;
    END
  END EXT_RDATABUS[7]
  PIN EXT_RDATABUS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 387.835000 0.070000 387.905000 ;
    END
  END EXT_RDATABUS[6]
  PIN EXT_RDATABUS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 394.835000 0.070000 394.905000 ;
    END
  END EXT_RDATABUS[5]
  PIN EXT_RDATABUS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 401.835000 0.070000 401.905000 ;
    END
  END EXT_RDATABUS[4]
  PIN EXT_RDATABUS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 408.835000 0.070000 408.905000 ;
    END
  END EXT_RDATABUS[3]
  PIN EXT_RDATABUS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 415.835000 0.070000 415.905000 ;
    END
  END EXT_RDATABUS[2]
  PIN EXT_RDATABUS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 422.835000 0.070000 422.905000 ;
    END
  END EXT_RDATABUS[1]
  PIN EXT_RDATABUS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 429.835000 0.070000 429.905000 ;
    END
  END EXT_RDATABUS[0]
  PIN EXT_WDATABUS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 411.915000 649.990000 411.985000 ;
    END
  END EXT_WDATABUS[31]
  PIN EXT_WDATABUS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 406.315000 649.990000 406.385000 ;
    END
  END EXT_WDATABUS[30]
  PIN EXT_WDATABUS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 400.715000 649.990000 400.785000 ;
    END
  END EXT_WDATABUS[29]
  PIN EXT_WDATABUS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 395.115000 649.990000 395.185000 ;
    END
  END EXT_WDATABUS[28]
  PIN EXT_WDATABUS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 389.515000 649.990000 389.585000 ;
    END
  END EXT_WDATABUS[27]
  PIN EXT_WDATABUS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 383.915000 649.990000 383.985000 ;
    END
  END EXT_WDATABUS[26]
  PIN EXT_WDATABUS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 378.315000 649.990000 378.385000 ;
    END
  END EXT_WDATABUS[25]
  PIN EXT_WDATABUS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 372.715000 649.990000 372.785000 ;
    END
  END EXT_WDATABUS[24]
  PIN EXT_WDATABUS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 367.115000 649.990000 367.185000 ;
    END
  END EXT_WDATABUS[23]
  PIN EXT_WDATABUS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 361.515000 649.990000 361.585000 ;
    END
  END EXT_WDATABUS[22]
  PIN EXT_WDATABUS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 355.915000 649.990000 355.985000 ;
    END
  END EXT_WDATABUS[21]
  PIN EXT_WDATABUS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 350.315000 649.990000 350.385000 ;
    END
  END EXT_WDATABUS[20]
  PIN EXT_WDATABUS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 344.715000 649.990000 344.785000 ;
    END
  END EXT_WDATABUS[19]
  PIN EXT_WDATABUS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 339.115000 649.990000 339.185000 ;
    END
  END EXT_WDATABUS[18]
  PIN EXT_WDATABUS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 333.515000 649.990000 333.585000 ;
    END
  END EXT_WDATABUS[17]
  PIN EXT_WDATABUS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 327.915000 649.990000 327.985000 ;
    END
  END EXT_WDATABUS[16]
  PIN EXT_WDATABUS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 322.315000 649.990000 322.385000 ;
    END
  END EXT_WDATABUS[15]
  PIN EXT_WDATABUS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 316.715000 649.990000 316.785000 ;
    END
  END EXT_WDATABUS[14]
  PIN EXT_WDATABUS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 311.115000 649.990000 311.185000 ;
    END
  END EXT_WDATABUS[13]
  PIN EXT_WDATABUS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 305.515000 649.990000 305.585000 ;
    END
  END EXT_WDATABUS[12]
  PIN EXT_WDATABUS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 299.915000 649.990000 299.985000 ;
    END
  END EXT_WDATABUS[11]
  PIN EXT_WDATABUS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 294.315000 649.990000 294.385000 ;
    END
  END EXT_WDATABUS[10]
  PIN EXT_WDATABUS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 288.715000 649.990000 288.785000 ;
    END
  END EXT_WDATABUS[9]
  PIN EXT_WDATABUS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 283.115000 649.990000 283.185000 ;
    END
  END EXT_WDATABUS[8]
  PIN EXT_WDATABUS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 277.515000 649.990000 277.585000 ;
    END
  END EXT_WDATABUS[7]
  PIN EXT_WDATABUS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 271.915000 649.990000 271.985000 ;
    END
  END EXT_WDATABUS[6]
  PIN EXT_WDATABUS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 266.315000 649.990000 266.385000 ;
    END
  END EXT_WDATABUS[5]
  PIN EXT_WDATABUS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 260.715000 649.990000 260.785000 ;
    END
  END EXT_WDATABUS[4]
  PIN EXT_WDATABUS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 255.115000 649.990000 255.185000 ;
    END
  END EXT_WDATABUS[3]
  PIN EXT_WDATABUS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 249.515000 649.990000 249.585000 ;
    END
  END EXT_WDATABUS[2]
  PIN EXT_WDATABUS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 243.915000 649.990000 243.985000 ;
    END
  END EXT_WDATABUS[1]
  PIN EXT_WDATABUS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 649.920000 238.315000 649.990000 238.385000 ;
    END
  END EXT_WDATABUS[0]
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 649.990000 650.020000 ;
    LAYER metal2 ;
      RECT 457.910000 649.880000 649.990000 650.020000 ;
      RECT 450.310000 649.880000 457.700000 650.020000 ;
      RECT 442.710000 649.880000 450.100000 650.020000 ;
      RECT 435.110000 649.880000 442.500000 650.020000 ;
      RECT 427.510000 649.880000 434.900000 650.020000 ;
      RECT 419.910000 649.880000 427.300000 650.020000 ;
      RECT 412.310000 649.880000 419.700000 650.020000 ;
      RECT 404.710000 649.880000 412.100000 650.020000 ;
      RECT 397.110000 649.880000 404.500000 650.020000 ;
      RECT 389.510000 649.880000 396.900000 650.020000 ;
      RECT 381.910000 649.880000 389.300000 650.020000 ;
      RECT 374.310000 649.880000 381.700000 650.020000 ;
      RECT 366.710000 649.880000 374.100000 650.020000 ;
      RECT 359.110000 649.880000 366.500000 650.020000 ;
      RECT 351.510000 649.880000 358.900000 650.020000 ;
      RECT 343.910000 649.880000 351.300000 650.020000 ;
      RECT 336.310000 649.880000 343.700000 650.020000 ;
      RECT 328.710000 649.880000 336.100000 650.020000 ;
      RECT 321.110000 649.880000 328.500000 650.020000 ;
      RECT 313.510000 649.880000 320.900000 650.020000 ;
      RECT 305.910000 649.880000 313.300000 650.020000 ;
      RECT 298.310000 649.880000 305.700000 650.020000 ;
      RECT 290.710000 649.880000 298.100000 650.020000 ;
      RECT 283.110000 649.880000 290.500000 650.020000 ;
      RECT 275.510000 649.880000 282.900000 650.020000 ;
      RECT 267.910000 649.880000 275.300000 650.020000 ;
      RECT 260.310000 649.880000 267.700000 650.020000 ;
      RECT 252.710000 649.880000 260.100000 650.020000 ;
      RECT 245.110000 649.880000 252.500000 650.020000 ;
      RECT 237.510000 649.880000 244.900000 650.020000 ;
      RECT 229.910000 649.880000 237.300000 650.020000 ;
      RECT 222.310000 649.880000 229.700000 650.020000 ;
      RECT 214.710000 649.880000 222.100000 650.020000 ;
      RECT 207.110000 649.880000 214.500000 650.020000 ;
      RECT 199.510000 649.880000 206.900000 650.020000 ;
      RECT 191.910000 649.880000 199.300000 650.020000 ;
      RECT 0.000000 649.880000 191.700000 650.020000 ;
      RECT 0.000000 436.975000 649.990000 649.880000 ;
      RECT 0.140000 436.765000 649.990000 436.975000 ;
      RECT 0.000000 429.975000 649.990000 436.765000 ;
      RECT 0.140000 429.765000 649.990000 429.975000 ;
      RECT 0.000000 422.975000 649.990000 429.765000 ;
      RECT 0.140000 422.765000 649.990000 422.975000 ;
      RECT 0.000000 415.975000 649.990000 422.765000 ;
      RECT 0.140000 415.765000 649.990000 415.975000 ;
      RECT 0.000000 412.055000 649.990000 415.765000 ;
      RECT 0.000000 411.845000 649.850000 412.055000 ;
      RECT 0.000000 408.975000 649.990000 411.845000 ;
      RECT 0.140000 408.765000 649.990000 408.975000 ;
      RECT 0.000000 406.455000 649.990000 408.765000 ;
      RECT 0.000000 406.245000 649.850000 406.455000 ;
      RECT 0.000000 401.975000 649.990000 406.245000 ;
      RECT 0.140000 401.765000 649.990000 401.975000 ;
      RECT 0.000000 400.855000 649.990000 401.765000 ;
      RECT 0.000000 400.645000 649.850000 400.855000 ;
      RECT 0.000000 395.255000 649.990000 400.645000 ;
      RECT 0.000000 395.045000 649.850000 395.255000 ;
      RECT 0.000000 394.975000 649.990000 395.045000 ;
      RECT 0.140000 394.765000 649.990000 394.975000 ;
      RECT 0.000000 389.655000 649.990000 394.765000 ;
      RECT 0.000000 389.445000 649.850000 389.655000 ;
      RECT 0.000000 387.975000 649.990000 389.445000 ;
      RECT 0.140000 387.765000 649.990000 387.975000 ;
      RECT 0.000000 384.055000 649.990000 387.765000 ;
      RECT 0.000000 383.845000 649.850000 384.055000 ;
      RECT 0.000000 380.975000 649.990000 383.845000 ;
      RECT 0.140000 380.765000 649.990000 380.975000 ;
      RECT 0.000000 378.455000 649.990000 380.765000 ;
      RECT 0.000000 378.245000 649.850000 378.455000 ;
      RECT 0.000000 373.975000 649.990000 378.245000 ;
      RECT 0.140000 373.765000 649.990000 373.975000 ;
      RECT 0.000000 372.855000 649.990000 373.765000 ;
      RECT 0.000000 372.645000 649.850000 372.855000 ;
      RECT 0.000000 367.255000 649.990000 372.645000 ;
      RECT 0.000000 367.045000 649.850000 367.255000 ;
      RECT 0.000000 366.975000 649.990000 367.045000 ;
      RECT 0.140000 366.765000 649.990000 366.975000 ;
      RECT 0.000000 361.655000 649.990000 366.765000 ;
      RECT 0.000000 361.445000 649.850000 361.655000 ;
      RECT 0.000000 359.975000 649.990000 361.445000 ;
      RECT 0.140000 359.765000 649.990000 359.975000 ;
      RECT 0.000000 356.055000 649.990000 359.765000 ;
      RECT 0.000000 355.845000 649.850000 356.055000 ;
      RECT 0.000000 352.975000 649.990000 355.845000 ;
      RECT 0.140000 352.765000 649.990000 352.975000 ;
      RECT 0.000000 350.455000 649.990000 352.765000 ;
      RECT 0.000000 350.245000 649.850000 350.455000 ;
      RECT 0.000000 345.975000 649.990000 350.245000 ;
      RECT 0.140000 345.765000 649.990000 345.975000 ;
      RECT 0.000000 344.855000 649.990000 345.765000 ;
      RECT 0.000000 344.645000 649.850000 344.855000 ;
      RECT 0.000000 339.255000 649.990000 344.645000 ;
      RECT 0.000000 339.045000 649.850000 339.255000 ;
      RECT 0.000000 338.975000 649.990000 339.045000 ;
      RECT 0.140000 338.765000 649.990000 338.975000 ;
      RECT 0.000000 333.655000 649.990000 338.765000 ;
      RECT 0.000000 333.445000 649.850000 333.655000 ;
      RECT 0.000000 331.975000 649.990000 333.445000 ;
      RECT 0.140000 331.765000 649.990000 331.975000 ;
      RECT 0.000000 328.055000 649.990000 331.765000 ;
      RECT 0.000000 327.845000 649.850000 328.055000 ;
      RECT 0.000000 324.975000 649.990000 327.845000 ;
      RECT 0.140000 324.765000 649.990000 324.975000 ;
      RECT 0.000000 322.455000 649.990000 324.765000 ;
      RECT 0.000000 322.245000 649.850000 322.455000 ;
      RECT 0.000000 317.975000 649.990000 322.245000 ;
      RECT 0.140000 317.765000 649.990000 317.975000 ;
      RECT 0.000000 316.855000 649.990000 317.765000 ;
      RECT 0.000000 316.645000 649.850000 316.855000 ;
      RECT 0.000000 311.255000 649.990000 316.645000 ;
      RECT 0.000000 311.045000 649.850000 311.255000 ;
      RECT 0.000000 310.975000 649.990000 311.045000 ;
      RECT 0.140000 310.765000 649.990000 310.975000 ;
      RECT 0.000000 305.655000 649.990000 310.765000 ;
      RECT 0.000000 305.445000 649.850000 305.655000 ;
      RECT 0.000000 303.975000 649.990000 305.445000 ;
      RECT 0.140000 303.765000 649.990000 303.975000 ;
      RECT 0.000000 300.055000 649.990000 303.765000 ;
      RECT 0.000000 299.845000 649.850000 300.055000 ;
      RECT 0.000000 296.975000 649.990000 299.845000 ;
      RECT 0.140000 296.765000 649.990000 296.975000 ;
      RECT 0.000000 294.455000 649.990000 296.765000 ;
      RECT 0.000000 294.245000 649.850000 294.455000 ;
      RECT 0.000000 289.975000 649.990000 294.245000 ;
      RECT 0.140000 289.765000 649.990000 289.975000 ;
      RECT 0.000000 288.855000 649.990000 289.765000 ;
      RECT 0.000000 288.645000 649.850000 288.855000 ;
      RECT 0.000000 283.255000 649.990000 288.645000 ;
      RECT 0.000000 283.045000 649.850000 283.255000 ;
      RECT 0.000000 282.975000 649.990000 283.045000 ;
      RECT 0.140000 282.765000 649.990000 282.975000 ;
      RECT 0.000000 277.655000 649.990000 282.765000 ;
      RECT 0.000000 277.445000 649.850000 277.655000 ;
      RECT 0.000000 275.975000 649.990000 277.445000 ;
      RECT 0.140000 275.765000 649.990000 275.975000 ;
      RECT 0.000000 272.055000 649.990000 275.765000 ;
      RECT 0.000000 271.845000 649.850000 272.055000 ;
      RECT 0.000000 268.975000 649.990000 271.845000 ;
      RECT 0.140000 268.765000 649.990000 268.975000 ;
      RECT 0.000000 266.455000 649.990000 268.765000 ;
      RECT 0.000000 266.245000 649.850000 266.455000 ;
      RECT 0.000000 261.975000 649.990000 266.245000 ;
      RECT 0.140000 261.765000 649.990000 261.975000 ;
      RECT 0.000000 260.855000 649.990000 261.765000 ;
      RECT 0.000000 260.645000 649.850000 260.855000 ;
      RECT 0.000000 255.255000 649.990000 260.645000 ;
      RECT 0.000000 255.045000 649.850000 255.255000 ;
      RECT 0.000000 254.975000 649.990000 255.045000 ;
      RECT 0.140000 254.765000 649.990000 254.975000 ;
      RECT 0.000000 249.655000 649.990000 254.765000 ;
      RECT 0.000000 249.445000 649.850000 249.655000 ;
      RECT 0.000000 247.975000 649.990000 249.445000 ;
      RECT 0.140000 247.765000 649.990000 247.975000 ;
      RECT 0.000000 244.055000 649.990000 247.765000 ;
      RECT 0.000000 243.845000 649.850000 244.055000 ;
      RECT 0.000000 240.975000 649.990000 243.845000 ;
      RECT 0.140000 240.765000 649.990000 240.975000 ;
      RECT 0.000000 238.455000 649.990000 240.765000 ;
      RECT 0.000000 238.245000 649.850000 238.455000 ;
      RECT 0.000000 233.975000 649.990000 238.245000 ;
      RECT 0.140000 233.765000 649.990000 233.975000 ;
      RECT 0.000000 226.975000 649.990000 233.765000 ;
      RECT 0.140000 226.765000 649.990000 226.975000 ;
      RECT 0.000000 219.975000 649.990000 226.765000 ;
      RECT 0.140000 219.765000 649.990000 219.975000 ;
      RECT 0.000000 212.975000 649.990000 219.765000 ;
      RECT 0.140000 212.765000 649.990000 212.975000 ;
      RECT 0.000000 0.000000 649.990000 212.765000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 649.990000 650.020000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 649.990000 650.020000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 649.990000 650.020000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 649.990000 650.020000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 649.990000 650.020000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 649.990000 650.020000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 649.990000 650.020000 ;
    LAYER metal10 ;
      RECT 0.000000 0.000000 649.990000 650.020000 ;
  END
END ensc450

END LIBRARY
