/local-scratch/localhome/escmc38/Desktop/ensc450/project/ensc450_system/BE_045/inputs/SRAM.lef