##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Sat Apr 17 14:47:07 2021
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core_adapter
  CLASS BLOCK ;
  SIZE 259.920000 BY 259.980000 ;
  FOREIGN core_adapter 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
  END clk
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.780000 259.910000 35.850000 259.980000 ;
    END
  END resetn
  PIN addr_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.630000 259.910000 38.700000 259.980000 ;
    END
  END addr_in[31]
  PIN addr_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.480000 259.910000 41.550000 259.980000 ;
    END
  END addr_in[30]
  PIN addr_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 44.330000 259.910000 44.400000 259.980000 ;
    END
  END addr_in[29]
  PIN addr_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 47.180000 259.910000 47.250000 259.980000 ;
    END
  END addr_in[28]
  PIN addr_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.030000 259.910000 50.100000 259.980000 ;
    END
  END addr_in[27]
  PIN addr_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.880000 259.910000 52.950000 259.980000 ;
    END
  END addr_in[26]
  PIN addr_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 55.730000 259.910000 55.800000 259.980000 ;
    END
  END addr_in[25]
  PIN addr_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.580000 259.910000 58.650000 259.980000 ;
    END
  END addr_in[24]
  PIN addr_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 61.430000 259.910000 61.500000 259.980000 ;
    END
  END addr_in[23]
  PIN addr_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.280000 259.910000 64.350000 259.980000 ;
    END
  END addr_in[22]
  PIN addr_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.130000 259.910000 67.200000 259.980000 ;
    END
  END addr_in[21]
  PIN addr_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.980000 259.910000 70.050000 259.980000 ;
    END
  END addr_in[20]
  PIN addr_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 72.830000 259.910000 72.900000 259.980000 ;
    END
  END addr_in[19]
  PIN addr_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 75.680000 259.910000 75.750000 259.980000 ;
    END
  END addr_in[18]
  PIN addr_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 78.530000 259.910000 78.600000 259.980000 ;
    END
  END addr_in[17]
  PIN addr_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.380000 259.910000 81.450000 259.980000 ;
    END
  END addr_in[16]
  PIN addr_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.230000 259.910000 84.300000 259.980000 ;
    END
  END addr_in[15]
  PIN addr_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 87.080000 259.910000 87.150000 259.980000 ;
    END
  END addr_in[14]
  PIN addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 89.930000 259.910000 90.000000 259.980000 ;
    END
  END addr_in[13]
  PIN addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.780000 259.910000 92.850000 259.980000 ;
    END
  END addr_in[12]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 95.630000 259.910000 95.700000 259.980000 ;
    END
  END addr_in[11]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.480000 259.910000 98.550000 259.980000 ;
    END
  END addr_in[10]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.330000 259.910000 101.400000 259.980000 ;
    END
  END addr_in[9]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 104.180000 259.910000 104.250000 259.980000 ;
    END
  END addr_in[8]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.030000 259.910000 107.100000 259.980000 ;
    END
  END addr_in[7]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 109.880000 259.910000 109.950000 259.980000 ;
    END
  END addr_in[6]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 112.730000 259.910000 112.800000 259.980000 ;
    END
  END addr_in[5]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 115.580000 259.910000 115.650000 259.980000 ;
    END
  END addr_in[4]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 118.430000 259.910000 118.500000 259.980000 ;
    END
  END addr_in[3]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.280000 259.910000 121.350000 259.980000 ;
    END
  END addr_in[2]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 124.130000 259.910000 124.200000 259.980000 ;
    END
  END addr_in[1]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 126.980000 259.910000 127.050000 259.980000 ;
    END
  END addr_in[0]
  PIN mr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 129.830000 259.910000 129.900000 259.980000 ;
    END
  END mr
  PIN mw
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 132.680000 259.910000 132.750000 259.980000 ;
    END
  END mw
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 135.530000 259.910000 135.600000 259.980000 ;
    END
  END data_in[31]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 138.380000 259.910000 138.450000 259.980000 ;
    END
  END data_in[30]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 141.230000 259.910000 141.300000 259.980000 ;
    END
  END data_in[29]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 144.080000 259.910000 144.150000 259.980000 ;
    END
  END data_in[28]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 146.930000 259.910000 147.000000 259.980000 ;
    END
  END data_in[27]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 149.780000 259.910000 149.850000 259.980000 ;
    END
  END data_in[26]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 152.630000 259.910000 152.700000 259.980000 ;
    END
  END data_in[25]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 155.480000 259.910000 155.550000 259.980000 ;
    END
  END data_in[24]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 158.330000 259.910000 158.400000 259.980000 ;
    END
  END data_in[23]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 161.180000 259.910000 161.250000 259.980000 ;
    END
  END data_in[22]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 164.030000 259.910000 164.100000 259.980000 ;
    END
  END data_in[21]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 166.880000 259.910000 166.950000 259.980000 ;
    END
  END data_in[20]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 169.730000 259.910000 169.800000 259.980000 ;
    END
  END data_in[19]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 172.580000 259.910000 172.650000 259.980000 ;
    END
  END data_in[18]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 175.430000 259.910000 175.500000 259.980000 ;
    END
  END data_in[17]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 178.280000 259.910000 178.350000 259.980000 ;
    END
  END data_in[16]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 181.130000 259.910000 181.200000 259.980000 ;
    END
  END data_in[15]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 183.980000 259.910000 184.050000 259.980000 ;
    END
  END data_in[14]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 186.830000 259.910000 186.900000 259.980000 ;
    END
  END data_in[13]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 189.680000 259.910000 189.750000 259.980000 ;
    END
  END data_in[12]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 192.530000 259.910000 192.600000 259.980000 ;
    END
  END data_in[11]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 195.380000 259.910000 195.450000 259.980000 ;
    END
  END data_in[10]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 198.230000 259.910000 198.300000 259.980000 ;
    END
  END data_in[9]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 201.080000 259.910000 201.150000 259.980000 ;
    END
  END data_in[8]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 203.930000 259.910000 204.000000 259.980000 ;
    END
  END data_in[7]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 206.780000 259.910000 206.850000 259.980000 ;
    END
  END data_in[6]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 209.630000 259.910000 209.700000 259.980000 ;
    END
  END data_in[5]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 212.480000 259.910000 212.550000 259.980000 ;
    END
  END data_in[4]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 215.330000 259.910000 215.400000 259.980000 ;
    END
  END data_in[3]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 218.180000 259.910000 218.250000 259.980000 ;
    END
  END data_in[2]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 221.030000 259.910000 221.100000 259.980000 ;
    END
  END data_in[1]
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 223.880000 259.910000 223.950000 259.980000 ;
    END
  END data_in[0]
  PIN data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 73.815000 0.070000 73.885000 ;
    END
  END data_out[31]
  PIN data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 77.315000 0.070000 77.385000 ;
    END
  END data_out[30]
  PIN data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 80.815000 0.070000 80.885000 ;
    END
  END data_out[29]
  PIN data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 84.315000 0.070000 84.385000 ;
    END
  END data_out[28]
  PIN data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 87.815000 0.070000 87.885000 ;
    END
  END data_out[27]
  PIN data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 91.315000 0.070000 91.385000 ;
    END
  END data_out[26]
  PIN data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 94.815000 0.070000 94.885000 ;
    END
  END data_out[25]
  PIN data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 98.315000 0.070000 98.385000 ;
    END
  END data_out[24]
  PIN data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 101.815000 0.070000 101.885000 ;
    END
  END data_out[23]
  PIN data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 105.315000 0.070000 105.385000 ;
    END
  END data_out[22]
  PIN data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 108.815000 0.070000 108.885000 ;
    END
  END data_out[21]
  PIN data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 112.315000 0.070000 112.385000 ;
    END
  END data_out[20]
  PIN data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 115.815000 0.070000 115.885000 ;
    END
  END data_out[19]
  PIN data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 119.315000 0.070000 119.385000 ;
    END
  END data_out[18]
  PIN data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 122.815000 0.070000 122.885000 ;
    END
  END data_out[17]
  PIN data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 126.315000 0.070000 126.385000 ;
    END
  END data_out[16]
  PIN data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 129.815000 0.070000 129.885000 ;
    END
  END data_out[15]
  PIN data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 133.315000 0.070000 133.385000 ;
    END
  END data_out[14]
  PIN data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 136.815000 0.070000 136.885000 ;
    END
  END data_out[13]
  PIN data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 140.315000 0.070000 140.385000 ;
    END
  END data_out[12]
  PIN data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 143.815000 0.070000 143.885000 ;
    END
  END data_out[11]
  PIN data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 147.315000 0.070000 147.385000 ;
    END
  END data_out[10]
  PIN data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 150.815000 0.070000 150.885000 ;
    END
  END data_out[9]
  PIN data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 154.315000 0.070000 154.385000 ;
    END
  END data_out[8]
  PIN data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 157.815000 0.070000 157.885000 ;
    END
  END data_out[7]
  PIN data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 161.315000 0.070000 161.385000 ;
    END
  END data_out[6]
  PIN data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 164.815000 0.070000 164.885000 ;
    END
  END data_out[5]
  PIN data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 168.315000 0.070000 168.385000 ;
    END
  END data_out[4]
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 171.815000 0.070000 171.885000 ;
    END
  END data_out[3]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 175.315000 0.070000 175.385000 ;
    END
  END data_out[2]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 178.815000 0.070000 178.885000 ;
    END
  END data_out[1]
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 182.315000 0.070000 182.385000 ;
    END
  END data_out[0]
  PIN nready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.000000 185.815000 0.070000 185.885000 ;
    END
  END nready
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 259.920000 259.980000 ;
    LAYER metal2 ;
      RECT 224.020000 259.840000 259.920000 259.980000 ;
      RECT 221.170000 259.840000 223.810000 259.980000 ;
      RECT 218.320000 259.840000 220.960000 259.980000 ;
      RECT 215.470000 259.840000 218.110000 259.980000 ;
      RECT 212.620000 259.840000 215.260000 259.980000 ;
      RECT 209.770000 259.840000 212.410000 259.980000 ;
      RECT 206.920000 259.840000 209.560000 259.980000 ;
      RECT 204.070000 259.840000 206.710000 259.980000 ;
      RECT 201.220000 259.840000 203.860000 259.980000 ;
      RECT 198.370000 259.840000 201.010000 259.980000 ;
      RECT 195.520000 259.840000 198.160000 259.980000 ;
      RECT 192.670000 259.840000 195.310000 259.980000 ;
      RECT 189.820000 259.840000 192.460000 259.980000 ;
      RECT 186.970000 259.840000 189.610000 259.980000 ;
      RECT 184.120000 259.840000 186.760000 259.980000 ;
      RECT 181.270000 259.840000 183.910000 259.980000 ;
      RECT 178.420000 259.840000 181.060000 259.980000 ;
      RECT 175.570000 259.840000 178.210000 259.980000 ;
      RECT 172.720000 259.840000 175.360000 259.980000 ;
      RECT 169.870000 259.840000 172.510000 259.980000 ;
      RECT 167.020000 259.840000 169.660000 259.980000 ;
      RECT 164.170000 259.840000 166.810000 259.980000 ;
      RECT 161.320000 259.840000 163.960000 259.980000 ;
      RECT 158.470000 259.840000 161.110000 259.980000 ;
      RECT 155.620000 259.840000 158.260000 259.980000 ;
      RECT 152.770000 259.840000 155.410000 259.980000 ;
      RECT 149.920000 259.840000 152.560000 259.980000 ;
      RECT 147.070000 259.840000 149.710000 259.980000 ;
      RECT 144.220000 259.840000 146.860000 259.980000 ;
      RECT 141.370000 259.840000 144.010000 259.980000 ;
      RECT 138.520000 259.840000 141.160000 259.980000 ;
      RECT 135.670000 259.840000 138.310000 259.980000 ;
      RECT 132.820000 259.840000 135.460000 259.980000 ;
      RECT 129.970000 259.840000 132.610000 259.980000 ;
      RECT 127.120000 259.840000 129.760000 259.980000 ;
      RECT 124.270000 259.840000 126.910000 259.980000 ;
      RECT 121.420000 259.840000 124.060000 259.980000 ;
      RECT 118.570000 259.840000 121.210000 259.980000 ;
      RECT 115.720000 259.840000 118.360000 259.980000 ;
      RECT 112.870000 259.840000 115.510000 259.980000 ;
      RECT 110.020000 259.840000 112.660000 259.980000 ;
      RECT 107.170000 259.840000 109.810000 259.980000 ;
      RECT 104.320000 259.840000 106.960000 259.980000 ;
      RECT 101.470000 259.840000 104.110000 259.980000 ;
      RECT 98.620000 259.840000 101.260000 259.980000 ;
      RECT 95.770000 259.840000 98.410000 259.980000 ;
      RECT 92.920000 259.840000 95.560000 259.980000 ;
      RECT 90.070000 259.840000 92.710000 259.980000 ;
      RECT 87.220000 259.840000 89.860000 259.980000 ;
      RECT 84.370000 259.840000 87.010000 259.980000 ;
      RECT 81.520000 259.840000 84.160000 259.980000 ;
      RECT 78.670000 259.840000 81.310000 259.980000 ;
      RECT 75.820000 259.840000 78.460000 259.980000 ;
      RECT 72.970000 259.840000 75.610000 259.980000 ;
      RECT 70.120000 259.840000 72.760000 259.980000 ;
      RECT 67.270000 259.840000 69.910000 259.980000 ;
      RECT 64.420000 259.840000 67.060000 259.980000 ;
      RECT 61.570000 259.840000 64.210000 259.980000 ;
      RECT 58.720000 259.840000 61.360000 259.980000 ;
      RECT 55.870000 259.840000 58.510000 259.980000 ;
      RECT 53.020000 259.840000 55.660000 259.980000 ;
      RECT 50.170000 259.840000 52.810000 259.980000 ;
      RECT 47.320000 259.840000 49.960000 259.980000 ;
      RECT 44.470000 259.840000 47.110000 259.980000 ;
      RECT 41.620000 259.840000 44.260000 259.980000 ;
      RECT 38.770000 259.840000 41.410000 259.980000 ;
      RECT 35.920000 259.840000 38.560000 259.980000 ;
      RECT 0.000000 259.840000 35.710000 259.980000 ;
      RECT 0.000000 185.955000 259.920000 259.840000 ;
      RECT 0.140000 185.745000 259.920000 185.955000 ;
      RECT 0.000000 182.455000 259.920000 185.745000 ;
      RECT 0.140000 182.245000 259.920000 182.455000 ;
      RECT 0.000000 178.955000 259.920000 182.245000 ;
      RECT 0.140000 178.745000 259.920000 178.955000 ;
      RECT 0.000000 175.455000 259.920000 178.745000 ;
      RECT 0.140000 175.245000 259.920000 175.455000 ;
      RECT 0.000000 171.955000 259.920000 175.245000 ;
      RECT 0.140000 171.745000 259.920000 171.955000 ;
      RECT 0.000000 168.455000 259.920000 171.745000 ;
      RECT 0.140000 168.245000 259.920000 168.455000 ;
      RECT 0.000000 164.955000 259.920000 168.245000 ;
      RECT 0.140000 164.745000 259.920000 164.955000 ;
      RECT 0.000000 161.455000 259.920000 164.745000 ;
      RECT 0.140000 161.245000 259.920000 161.455000 ;
      RECT 0.000000 157.955000 259.920000 161.245000 ;
      RECT 0.140000 157.745000 259.920000 157.955000 ;
      RECT 0.000000 154.455000 259.920000 157.745000 ;
      RECT 0.140000 154.245000 259.920000 154.455000 ;
      RECT 0.000000 150.955000 259.920000 154.245000 ;
      RECT 0.140000 150.745000 259.920000 150.955000 ;
      RECT 0.000000 147.455000 259.920000 150.745000 ;
      RECT 0.140000 147.245000 259.920000 147.455000 ;
      RECT 0.000000 143.955000 259.920000 147.245000 ;
      RECT 0.140000 143.745000 259.920000 143.955000 ;
      RECT 0.000000 140.455000 259.920000 143.745000 ;
      RECT 0.140000 140.245000 259.920000 140.455000 ;
      RECT 0.000000 136.955000 259.920000 140.245000 ;
      RECT 0.140000 136.745000 259.920000 136.955000 ;
      RECT 0.000000 133.455000 259.920000 136.745000 ;
      RECT 0.140000 133.245000 259.920000 133.455000 ;
      RECT 0.000000 129.955000 259.920000 133.245000 ;
      RECT 0.140000 129.745000 259.920000 129.955000 ;
      RECT 0.000000 126.455000 259.920000 129.745000 ;
      RECT 0.140000 126.245000 259.920000 126.455000 ;
      RECT 0.000000 122.955000 259.920000 126.245000 ;
      RECT 0.140000 122.745000 259.920000 122.955000 ;
      RECT 0.000000 119.455000 259.920000 122.745000 ;
      RECT 0.140000 119.245000 259.920000 119.455000 ;
      RECT 0.000000 115.955000 259.920000 119.245000 ;
      RECT 0.140000 115.745000 259.920000 115.955000 ;
      RECT 0.000000 112.455000 259.920000 115.745000 ;
      RECT 0.140000 112.245000 259.920000 112.455000 ;
      RECT 0.000000 108.955000 259.920000 112.245000 ;
      RECT 0.140000 108.745000 259.920000 108.955000 ;
      RECT 0.000000 105.455000 259.920000 108.745000 ;
      RECT 0.140000 105.245000 259.920000 105.455000 ;
      RECT 0.000000 101.955000 259.920000 105.245000 ;
      RECT 0.140000 101.745000 259.920000 101.955000 ;
      RECT 0.000000 98.455000 259.920000 101.745000 ;
      RECT 0.140000 98.245000 259.920000 98.455000 ;
      RECT 0.000000 94.955000 259.920000 98.245000 ;
      RECT 0.140000 94.745000 259.920000 94.955000 ;
      RECT 0.000000 91.455000 259.920000 94.745000 ;
      RECT 0.140000 91.245000 259.920000 91.455000 ;
      RECT 0.000000 87.955000 259.920000 91.245000 ;
      RECT 0.140000 87.745000 259.920000 87.955000 ;
      RECT 0.000000 84.455000 259.920000 87.745000 ;
      RECT 0.140000 84.245000 259.920000 84.455000 ;
      RECT 0.000000 80.955000 259.920000 84.245000 ;
      RECT 0.140000 80.745000 259.920000 80.955000 ;
      RECT 0.000000 77.455000 259.920000 80.745000 ;
      RECT 0.140000 77.245000 259.920000 77.455000 ;
      RECT 0.000000 73.955000 259.920000 77.245000 ;
      RECT 0.140000 73.745000 259.920000 73.955000 ;
      RECT 0.000000 0.000000 259.920000 73.745000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 259.920000 259.980000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 259.920000 259.980000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 259.920000 259.980000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 259.920000 259.980000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 259.920000 259.980000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 259.920000 259.980000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 259.920000 259.980000 ;
    LAYER metal10 ;
      RECT 0.000000 0.000000 259.920000 259.980000 ;
  END
END core_adapter

END LIBRARY
